module hello_world;
   initial begin
      $display("Hello, Verilog World!");
   end
endmodule
